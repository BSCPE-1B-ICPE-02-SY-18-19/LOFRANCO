CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 6 110 10
176 80 1534 813
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
110100626 0
0
6 Title:
5 Name:
0
0
0
10
2 +V
167 280 224 0 1 3
0 4
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5130 0 0
2
43529.7 0
0
7 Pulser~
4 93 306 0 10 12
0 17 18 3 19 0 0 5 5 6
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
391 0 0
2
43529.7 1
0
9 CC 7-Seg~
183 873 292 0 18 19
10 10 9 8 2 7 6 5 20 21
2 2 2 2 2 2 2 2 2
0
0 0 21104 0
6 BLUECC
-76 -3 -34 5
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3124 0 0
2
43529.7 2
0
9 2-In AND~
219 604 213 0 3 22
0 16 12 15
0
0 0 624 0
6 74LS08
-25 22 17 30
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3421 0 0
2
43529.7 3
0
9 2-In AND~
219 477 214 0 3 22
0 13 14 16
0
0 0 624 0
6 74LS08
-24 21 18 29
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
8157 0 0
2
43529.7 4
0
6 74112~
219 658 330 0 7 32
0 4 15 3 15 4 22 11
0
0 0 4720 0
5 74112
-72 -22 -37 -14
3 FFD
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
5572 0 0
2
43529.7 5
0
6 74112~
219 532 330 0 7 32
0 4 16 3 16 4 23 12
0
0 0 4720 0
5 74112
-72 -23 -37 -15
3 FFC
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
8901 0 0
2
43529.7 6
0
6 74112~
219 406 330 0 7 32
0 4 13 3 13 4 24 14
0
0 0 4720 0
5 74112
-71 -23 -36 -15
3 FFB
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
7361 0 0
2
43529.7 7
0
6 74112~
219 280 330 0 7 32
0 4 4 3 4 4 25 13
0
0 0 4720 0
5 74112
-72 -24 -37 -16
3 FFA
21 -62 42 -54
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
4747 0 0
2
43529.7 8
0
6 74LS48
188 774 403 0 14 29
0 11 12 14 13 26 27 5 6 7
2 8 9 10 28
0
0 0 4848 0
6 74LS48
-20 59 22 67
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
972 0 0
2
43529.7 9
0
35
10 4 2 0 0 8320 0 10 3 0 0 3
806 394
870 394
870 328
3 0 3 0 0 4096 0 9 0 0 10 2
250 303
250 359
2 1 4 0 0 4096 0 9 1 0 0 3
256 294
256 233
280 233
4 2 4 0 0 0 0 9 9 0 0 2
256 312
256 294
0 0 4 0 0 4096 0 0 0 6 13 2
326 267
326 342
1 1 4 0 0 4224 0 9 8 0 0 2
280 267
406 267
1 1 4 0 0 0 0 1 9 0 0 2
280 233
280 267
3 0 3 0 0 0 0 8 0 0 10 2
376 303
376 359
3 0 3 0 0 0 0 7 0 0 10 2
502 303
502 359
3 3 3 0 0 12416 0 2 6 0 0 5
117 297
169 297
169 359
628 359
628 303
5 5 4 0 0 128 0 7 6 0 0 2
532 342
658 342
5 5 4 0 0 0 0 8 7 0 0 2
406 342
532 342
5 5 4 0 0 0 0 9 8 0 0 2
280 342
406 342
7 7 5 0 0 4224 0 10 3 0 0 3
806 367
888 367
888 328
8 6 6 0 0 4224 0 10 3 0 0 3
806 376
882 376
882 328
9 5 7 0 0 4224 0 10 3 0 0 3
806 385
876 385
876 328
11 3 8 0 0 8320 0 10 3 0 0 3
806 403
864 403
864 328
12 2 9 0 0 8320 0 10 3 0 0 3
806 412
858 412
858 328
13 1 10 0 0 8320 0 10 3 0 0 3
806 421
852 421
852 328
1 7 11 0 0 8320 0 10 6 0 0 3
742 367
682 367
682 294
7 2 12 0 0 8320 0 7 10 0 0 3
556 294
556 376
742 376
7 4 13 0 0 8320 0 9 10 0 0 3
304 294
304 394
742 394
3 7 14 0 0 4224 0 10 8 0 0 3
742 385
430 385
430 294
2 3 15 0 0 4224 0 6 4 0 0 3
634 294
634 213
625 213
2 7 12 0 0 0 0 4 7 0 0 3
580 222
580 294
556 294
3 1 16 0 0 4096 0 5 4 0 0 4
498 214
567 214
567 204
580 204
2 3 16 0 0 4224 0 7 5 0 0 3
508 294
508 214
498 214
2 1 13 0 0 0 0 8 5 0 0 3
382 294
382 205
453 205
7 2 14 0 0 0 0 8 5 0 0 3
430 294
430 223
453 223
7 2 13 0 0 0 0 9 8 0 0 2
304 294
382 294
2 4 15 0 0 0 0 6 6 0 0 2
634 294
634 312
2 4 16 0 0 0 0 7 7 0 0 2
508 294
508 312
2 4 13 0 0 0 0 8 8 0 0 2
382 294
382 312
1 1 4 0 0 128 0 7 6 0 0 2
532 267
658 267
1 1 4 0 0 0 0 8 7 0 0 2
406 267
532 267
2
-21 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 37
27 13 582 48
36 20 572 43
37 LOFRANCO, JHON KENNETH C.		BSCPE - 1B
-32 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 35
228 97 916 153
239 105 904 141
35 BINARY 4-BIT SYNCHRONOUS UP COUNTER
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
